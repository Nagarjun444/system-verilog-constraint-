1)iam having 16bit of variable only single bit has to acess how to use of constraints
ex:4--->100
8---->1000
16---->10000
2)write a constraint to generate mul of 2 power?
3)write a constraint sunch that array size between 5 to 10 values of the array are in asscending/descending order ?
4)write a constraint to generate unique elements with out unique keyword?
5)how to delate/remove duplicate elements using queue?
6)how to delate/remove duplicate elements using associative array?
7)write a constraint to generate a variable with 0-31 bits should be 1,32-61 bits should be 0.
8)if we randomize a single bit variable for 10 times values should generate be like 101010101010.
9)we have a randomize variable with size of 32 bit data,but randomize only 12th bit.


//-----------D15------------------
1)generate odd number/even number ina fixed size array using $random
2)Write a constraint for 2D fixed size array randomization using Dynamic array ?
3)Write a constraint to generate the below pattern in dynamic array ?
0 1 0 2 0 3 0 4 0 5 0 
4)Pre Post Randomization examples
5)write a constraint to randmoly genrate 10 unquie numbers between 99 to 100
6)Write constraint to generate random values 25,27,30,36,40,45 without using "set membership". 
